magic
tech sky130B
magscale 1 2
timestamp 1667654173
<< metal4 >>
rect -2349 2039 2349 2080
rect -2349 -2039 2093 2039
rect 2329 -2039 2349 2039
rect -2349 -2080 2349 -2039
<< via4 >>
rect 2093 -2039 2329 2039
<< mimcap2 >>
rect -2269 1960 1731 2000
rect -2269 -1960 -2229 1960
rect 1691 -1960 1731 1960
rect -2269 -2000 1731 -1960
<< mimcap2contact >>
rect -2229 -1960 1691 1960
<< metal5 >>
rect 2051 2039 2371 2081
rect -2253 1960 1715 1984
rect -2253 -1960 -2229 1960
rect 1691 -1960 1715 1960
rect -2253 -1984 1715 -1960
rect 2051 -2039 2093 2039
rect 2329 -2039 2371 2039
rect 2051 -2081 2371 -2039
<< properties >>
string FIXED_BBOX -2349 -2080 1811 2080
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 20 l 20 val 815.2 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
